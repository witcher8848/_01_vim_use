module fifo (
    
);
begin
end
endmodule
